// The code is defined in the module which are similar to main functions in C language
// Here module is keyword
// andgate is module name
// The inputs and outputs are enclosed in the parenthesis
module andgate (a,b,y);

// defining inputs and outputs
input a,b;
output y;

// performing operation on the inputs and outputs and assigning the value to y
assign y = a&b;

// ending the module
endmodule

